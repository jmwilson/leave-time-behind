.SUBCKT LMERR_AMP PLUS MINUS OUT
R1 PLUS 0 1G
R2 MINUS 0 1G
R3 4 0 1G
D1 11 OUT _LMERR
.MODEL _LMERR D BV=1
V2 11 0 DC = 1.3
GB7 0 OUT VALUE {25E-6*V(9)}
EB9 3 0 VALUE {V(1)}
GB3 0 4 VALUE {1000*(V(PLUS,MINUS)-V(2))}
R5 3 9 1K
R7 0 2 10K
R8 2 1 300K
C4 4 0 10U
EB4 5 0 VALUE {V(4)}
R9 5 1 1
C5 1 0 .02U
D2 9 10 _D2_MOD
.MODEL _D2_MOD D BV=9
R10 OUT 0 48K
V5 10 0 DC = 5
.ENDS LMERR_AMP
